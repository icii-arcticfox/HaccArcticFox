module Settings;


/*[$^UseHardwareAcceleration true]*/
/*[$^RadiationValueWidth 32]*/
endmodule