module Settings;

//Switch to true when you want to use hardware acceleration
/*[$^UseHardwareAcceleration false]*/

//Don't change
/*[$^RadiationValueWidth 32]*/
endmodule