//[ExternalGroup RadiationReceiver]
/*[NormalChecks]*/
module HardwareAcceleratedHistogram(
);

//In this file you will implement you hardware accelerated histogram
endmodule