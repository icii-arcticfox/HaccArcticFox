module Settings;


/*[$^UseHardwareAcceleration false]*/
/*[$^RadiationValueWidth 32]*/

endmodule